import("EV3_common.cdl");

/*
 * MainTask:   主タスク       EV3 起動時から起動  優先度 EV3_MRUBY_VM_MAIN_PRIORITY
 */

//[domain(HRP2, "trusted")]
//[domain(HRP2, "nontrusted")]
region rDomainEV3 {
  /*----------- Main VM  -----------*/
	cell nMruby::tMruby MrubyMainVM {
		mrubyFile="$(MRUBY_LIB_DIR)/EV3_common.rb "
				"$(MRUBY_LIB_DIR)/RTOS.rb "
       			"$(MRUBY_LIB_DIR)/Speaker.rb "
				"$(MRUBY_LIB_DIR)/Button.rb "
				"$(MRUBY_LIB_DIR)/Motor.rb "
				"$(MRUBY_LIB_DIR)/UltrasonicSensor.rb "
				"$(MRUBY_LIB_DIR)/GyroSensor.rb "
				"$(MRUBY_LIB_DIR)/ColorSensor.rb "
				"$(MRUBY_LIB_DIR)/TouchSensor.rb "
				"$(MRUBY_LIB_DIR)/LED.rb "
				"$(MRUBY_LIB_DIR)/LCD.rb "
				"$(MRUBY_LIB_DIR)/Battery.rb "
				"$(MRUBY_LIB_DIR)/Balancer.rb "
        		"sharedmemory_def.rb "
        		"$(MRUBY_LIB_DIR)/SharedMemory.rb "
				"$(RUBY_FILE) "
				"$(APP_RB)";
		cInit = VM_TECSInitializer.eInitialize;
	};
	cell tTask MrubyMainTask {
	// 呼び口の結合 
		cBody = MrubyMainVM.eMrubyBody;
		//* 属性の設定
		taskAttribute = C_EXP("TA_ACT");
		priority = C_EXP("EV3_MRUBY_VM_MAIN_PRIORITY");
		systemStackSize = C_EXP("MRUBY_VM_STACK_SIZE");
	};

  /*-------*/
};


/*** Bridges ***/
generate( MrubyBridgePlugin, tTask, "" );
generate( MrubyBridgePlugin, tSemaphore, "" );

